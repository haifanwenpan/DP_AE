// CRC polynomial coefficients: x^32 + x^26 + x^23 + x^22 + x^16 + x^12 + x^11 + x^10 + x^8 + x^7 + x^5 + x^4 + x^2 + x + 1
//                              0x4C11DB7 (hex)
// CRC width:                   32 bits
// CRC shift direction:         left (big endian)
// Input word width:            144 bits
`default_nettype none
module CRC_32_DAT_144 (
    input  wire [ 31:0] CRC_IN,
    input  wire [143:0] DATA,
    output wire [ 31:0] CRC_OUT
);
  assign CRC_OUT[0] = CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[11] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[20] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[31] ^ DATA[0] ^ DATA[6] ^ DATA[9] ^ DATA[10] ^ DATA[12] ^ DATA[16] ^ DATA[24] ^ DATA[25] ^ DATA[26] ^ DATA[28] ^ DATA[29] ^ DATA[30] ^ DATA[31] ^ DATA[32] ^ DATA[34] ^ DATA[37] ^ DATA[44] ^ DATA[45] ^ DATA[47] ^ DATA[48] ^ DATA[50] ^ DATA[53] ^ DATA[54] ^ DATA[55] ^ DATA[58] ^ DATA[60] ^ DATA[61] ^ DATA[63] ^ DATA[65] ^ DATA[66] ^ DATA[67] ^ DATA[68] ^ DATA[72] ^ DATA[73] ^ DATA[79] ^ DATA[81] ^ DATA[82] ^ DATA[83] ^ DATA[84] ^ DATA[85] ^ DATA[87] ^ DATA[94] ^ DATA[95] ^ DATA[96] ^ DATA[97] ^ DATA[98] ^ DATA[99] ^ DATA[101] ^ DATA[103] ^ DATA[104] ^ DATA[106] ^ DATA[110] ^ DATA[111] ^ DATA[113] ^ DATA[114] ^ DATA[116] ^ DATA[117] ^ DATA[118] ^ DATA[119] ^ DATA[123] ^ DATA[125] ^ DATA[126] ^ DATA[127] ^ DATA[128] ^ DATA[132] ^ DATA[134] ^ DATA[135] ^ DATA[136] ^ DATA[137] ^ DATA[143];
  assign CRC_OUT[1] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[8] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[17] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[26] ^ CRC_IN[31] ^ DATA[0] ^ DATA[1] ^ DATA[6] ^ DATA[7] ^ DATA[9] ^ DATA[11] ^ DATA[12] ^ DATA[13] ^ DATA[16] ^ DATA[17] ^ DATA[24] ^ DATA[27] ^ DATA[28] ^ DATA[33] ^ DATA[34] ^ DATA[35] ^ DATA[37] ^ DATA[38] ^ DATA[44] ^ DATA[46] ^ DATA[47] ^ DATA[49] ^ DATA[50] ^ DATA[51] ^ DATA[53] ^ DATA[56] ^ DATA[58] ^ DATA[59] ^ DATA[60] ^ DATA[62] ^ DATA[63] ^ DATA[64] ^ DATA[65] ^ DATA[69] ^ DATA[72] ^ DATA[74] ^ DATA[79] ^ DATA[80] ^ DATA[81] ^ DATA[86] ^ DATA[87] ^ DATA[88] ^ DATA[94] ^ DATA[100] ^ DATA[101] ^ DATA[102] ^ DATA[103] ^ DATA[105] ^ DATA[106] ^ DATA[107] ^ DATA[110] ^ DATA[112] ^ DATA[113] ^ DATA[115] ^ DATA[116] ^ DATA[120] ^ DATA[123] ^ DATA[124] ^ DATA[125] ^ DATA[129] ^ DATA[132] ^ DATA[133] ^ DATA[134] ^ DATA[138] ^ DATA[143];
  assign CRC_OUT[2] = CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[9] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[18] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[27] ^ CRC_IN[31] ^ DATA[0] ^ DATA[1] ^ DATA[2] ^ DATA[6] ^ DATA[7] ^ DATA[8] ^ DATA[9] ^ DATA[13] ^ DATA[14] ^ DATA[16] ^ DATA[17] ^ DATA[18] ^ DATA[24] ^ DATA[26] ^ DATA[30] ^ DATA[31] ^ DATA[32] ^ DATA[35] ^ DATA[36] ^ DATA[37] ^ DATA[38] ^ DATA[39] ^ DATA[44] ^ DATA[51] ^ DATA[52] ^ DATA[53] ^ DATA[55] ^ DATA[57] ^ DATA[58] ^ DATA[59] ^ DATA[64] ^ DATA[67] ^ DATA[68] ^ DATA[70] ^ DATA[72] ^ DATA[75] ^ DATA[79] ^ DATA[80] ^ DATA[83] ^ DATA[84] ^ DATA[85] ^ DATA[88] ^ DATA[89] ^ DATA[94] ^ DATA[96] ^ DATA[97] ^ DATA[98] ^ DATA[99] ^ DATA[102] ^ DATA[107] ^ DATA[108] ^ DATA[110] ^ DATA[118] ^ DATA[119] ^ DATA[121] ^ DATA[123] ^ DATA[124] ^ DATA[127] ^ DATA[128] ^ DATA[130] ^ DATA[132] ^ DATA[133] ^ DATA[136] ^ DATA[137] ^ DATA[139] ^ DATA[143];
  assign CRC_OUT[3] = CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[19] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[28] ^ DATA[1] ^ DATA[2] ^ DATA[3] ^ DATA[7] ^ DATA[8] ^ DATA[9] ^ DATA[10] ^ DATA[14] ^ DATA[15] ^ DATA[17] ^ DATA[18] ^ DATA[19] ^ DATA[25] ^ DATA[27] ^ DATA[31] ^ DATA[32] ^ DATA[33] ^ DATA[36] ^ DATA[37] ^ DATA[38] ^ DATA[39] ^ DATA[40] ^ DATA[45] ^ DATA[52] ^ DATA[53] ^ DATA[54] ^ DATA[56] ^ DATA[58] ^ DATA[59] ^ DATA[60] ^ DATA[65] ^ DATA[68] ^ DATA[69] ^ DATA[71] ^ DATA[73] ^ DATA[76] ^ DATA[80] ^ DATA[81] ^ DATA[84] ^ DATA[85] ^ DATA[86] ^ DATA[89] ^ DATA[90] ^ DATA[95] ^ DATA[97] ^ DATA[98] ^ DATA[99] ^ DATA[100] ^ DATA[103] ^ DATA[108] ^ DATA[109] ^ DATA[111] ^ DATA[119] ^ DATA[120] ^ DATA[122] ^ DATA[124] ^ DATA[125] ^ DATA[128] ^ DATA[129] ^ DATA[131] ^ DATA[133] ^ DATA[134] ^ DATA[137] ^ DATA[138] ^ DATA[140];
  assign CRC_OUT[4] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[0] ^ DATA[2] ^ DATA[3] ^ DATA[4] ^ DATA[6] ^ DATA[8] ^ DATA[11] ^ DATA[12] ^ DATA[15] ^ DATA[18] ^ DATA[19] ^ DATA[20] ^ DATA[24] ^ DATA[25] ^ DATA[29] ^ DATA[30] ^ DATA[31] ^ DATA[33] ^ DATA[38] ^ DATA[39] ^ DATA[40] ^ DATA[41] ^ DATA[44] ^ DATA[45] ^ DATA[46] ^ DATA[47] ^ DATA[48] ^ DATA[50] ^ DATA[57] ^ DATA[58] ^ DATA[59] ^ DATA[63] ^ DATA[65] ^ DATA[67] ^ DATA[68] ^ DATA[69] ^ DATA[70] ^ DATA[73] ^ DATA[74] ^ DATA[77] ^ DATA[79] ^ DATA[83] ^ DATA[84] ^ DATA[86] ^ DATA[90] ^ DATA[91] ^ DATA[94] ^ DATA[95] ^ DATA[97] ^ DATA[100] ^ DATA[103] ^ DATA[106] ^ DATA[109] ^ DATA[111] ^ DATA[112] ^ DATA[113] ^ DATA[114] ^ DATA[116] ^ DATA[117] ^ DATA[118] ^ DATA[119] ^ DATA[120] ^ DATA[121] ^ DATA[127] ^ DATA[128] ^ DATA[129] ^ DATA[130] ^ DATA[136] ^ DATA[137] ^ DATA[138] ^ DATA[139] ^ DATA[141] ^ DATA[143];
  assign CRC_OUT[5] = CRC_IN[0] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[28] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[0] ^ DATA[1] ^ DATA[3] ^ DATA[4] ^ DATA[5] ^ DATA[6] ^ DATA[7] ^ DATA[10] ^ DATA[13] ^ DATA[19] ^ DATA[20] ^ DATA[21] ^ DATA[24] ^ DATA[28] ^ DATA[29] ^ DATA[37] ^ DATA[39] ^ DATA[40] ^ DATA[41] ^ DATA[42] ^ DATA[44] ^ DATA[46] ^ DATA[49] ^ DATA[50] ^ DATA[51] ^ DATA[53] ^ DATA[54] ^ DATA[55] ^ DATA[59] ^ DATA[61] ^ DATA[63] ^ DATA[64] ^ DATA[65] ^ DATA[67] ^ DATA[69] ^ DATA[70] ^ DATA[71] ^ DATA[72] ^ DATA[73] ^ DATA[74] ^ DATA[75] ^ DATA[78] ^ DATA[79] ^ DATA[80] ^ DATA[81] ^ DATA[82] ^ DATA[83] ^ DATA[91] ^ DATA[92] ^ DATA[94] ^ DATA[97] ^ DATA[99] ^ DATA[103] ^ DATA[106] ^ DATA[107] ^ DATA[111] ^ DATA[112] ^ DATA[115] ^ DATA[116] ^ DATA[120] ^ DATA[121] ^ DATA[122] ^ DATA[123] ^ DATA[125] ^ DATA[126] ^ DATA[127] ^ DATA[129] ^ DATA[130] ^ DATA[131] ^ DATA[132] ^ DATA[134] ^ DATA[135] ^ DATA[136] ^ DATA[138] ^ DATA[139] ^ DATA[140] ^ DATA[142] ^ DATA[143];
  assign CRC_OUT[6] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[27] ^ CRC_IN[28] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[1] ^ DATA[2] ^ DATA[4] ^ DATA[5] ^ DATA[6] ^ DATA[7] ^ DATA[8] ^ DATA[11] ^ DATA[14] ^ DATA[20] ^ DATA[21] ^ DATA[22] ^ DATA[25] ^ DATA[29] ^ DATA[30] ^ DATA[38] ^ DATA[40] ^ DATA[41] ^ DATA[42] ^ DATA[43] ^ DATA[45] ^ DATA[47] ^ DATA[50] ^ DATA[51] ^ DATA[52] ^ DATA[54] ^ DATA[55] ^ DATA[56] ^ DATA[60] ^ DATA[62] ^ DATA[64] ^ DATA[65] ^ DATA[66] ^ DATA[68] ^ DATA[70] ^ DATA[71] ^ DATA[72] ^ DATA[73] ^ DATA[74] ^ DATA[75] ^ DATA[76] ^ DATA[79] ^ DATA[80] ^ DATA[81] ^ DATA[82] ^ DATA[83] ^ DATA[84] ^ DATA[92] ^ DATA[93] ^ DATA[95] ^ DATA[98] ^ DATA[100] ^ DATA[104] ^ DATA[107] ^ DATA[108] ^ DATA[112] ^ DATA[113] ^ DATA[116] ^ DATA[117] ^ DATA[121] ^ DATA[122] ^ DATA[123] ^ DATA[124] ^ DATA[126] ^ DATA[127] ^ DATA[128] ^ DATA[130] ^ DATA[131] ^ DATA[132] ^ DATA[133] ^ DATA[135] ^ DATA[136] ^ DATA[137] ^ DATA[139] ^ DATA[140] ^ DATA[141] ^ DATA[143];
  assign CRC_OUT[7] = CRC_IN[4] ^ CRC_IN[7] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[14] ^ CRC_IN[17] ^ CRC_IN[19] ^ CRC_IN[21] ^ CRC_IN[23] ^ CRC_IN[26] ^ CRC_IN[28] ^ CRC_IN[29] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[0] ^ DATA[2] ^ DATA[3] ^ DATA[5] ^ DATA[7] ^ DATA[8] ^ DATA[10] ^ DATA[15] ^ DATA[16] ^ DATA[21] ^ DATA[22] ^ DATA[23] ^ DATA[24] ^ DATA[25] ^ DATA[28] ^ DATA[29] ^ DATA[32] ^ DATA[34] ^ DATA[37] ^ DATA[39] ^ DATA[41] ^ DATA[42] ^ DATA[43] ^ DATA[45] ^ DATA[46] ^ DATA[47] ^ DATA[50] ^ DATA[51] ^ DATA[52] ^ DATA[54] ^ DATA[56] ^ DATA[57] ^ DATA[58] ^ DATA[60] ^ DATA[68] ^ DATA[69] ^ DATA[71] ^ DATA[74] ^ DATA[75] ^ DATA[76] ^ DATA[77] ^ DATA[79] ^ DATA[80] ^ DATA[87] ^ DATA[93] ^ DATA[95] ^ DATA[97] ^ DATA[98] ^ DATA[103] ^ DATA[104] ^ DATA[105] ^ DATA[106] ^ DATA[108] ^ DATA[109] ^ DATA[110] ^ DATA[111] ^ DATA[116] ^ DATA[119] ^ DATA[122] ^ DATA[124] ^ DATA[126] ^ DATA[129] ^ DATA[131] ^ DATA[133] ^ DATA[135] ^ DATA[138] ^ DATA[140] ^ DATA[141] ^ DATA[142] ^ DATA[143];
  assign CRC_OUT[8] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[4] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[14] ^ CRC_IN[16] ^ CRC_IN[18] ^ CRC_IN[23] ^ CRC_IN[25] ^ CRC_IN[27] ^ CRC_IN[29] ^ CRC_IN[30] ^ DATA[0] ^ DATA[1] ^ DATA[3] ^ DATA[4] ^ DATA[8] ^ DATA[10] ^ DATA[11] ^ DATA[12] ^ DATA[17] ^ DATA[22] ^ DATA[23] ^ DATA[28] ^ DATA[31] ^ DATA[32] ^ DATA[33] ^ DATA[34] ^ DATA[35] ^ DATA[37] ^ DATA[38] ^ DATA[40] ^ DATA[42] ^ DATA[43] ^ DATA[45] ^ DATA[46] ^ DATA[50] ^ DATA[51] ^ DATA[52] ^ DATA[54] ^ DATA[57] ^ DATA[59] ^ DATA[60] ^ DATA[63] ^ DATA[65] ^ DATA[66] ^ DATA[67] ^ DATA[68] ^ DATA[69] ^ DATA[70] ^ DATA[73] ^ DATA[75] ^ DATA[76] ^ DATA[77] ^ DATA[78] ^ DATA[79] ^ DATA[80] ^ DATA[82] ^ DATA[83] ^ DATA[84] ^ DATA[85] ^ DATA[87] ^ DATA[88] ^ DATA[95] ^ DATA[97] ^ DATA[101] ^ DATA[103] ^ DATA[105] ^ DATA[107] ^ DATA[109] ^ DATA[112] ^ DATA[113] ^ DATA[114] ^ DATA[116] ^ DATA[118] ^ DATA[119] ^ DATA[120] ^ DATA[126] ^ DATA[128] ^ DATA[130] ^ DATA[135] ^ DATA[137] ^ DATA[139] ^ DATA[141] ^ DATA[142];
  assign CRC_OUT[9] = CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[5] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[15] ^ CRC_IN[17] ^ CRC_IN[19] ^ CRC_IN[24] ^ CRC_IN[26] ^ CRC_IN[28] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[1] ^ DATA[2] ^ DATA[4] ^ DATA[5] ^ DATA[9] ^ DATA[11] ^ DATA[12] ^ DATA[13] ^ DATA[18] ^ DATA[23] ^ DATA[24] ^ DATA[29] ^ DATA[32] ^ DATA[33] ^ DATA[34] ^ DATA[35] ^ DATA[36] ^ DATA[38] ^ DATA[39] ^ DATA[41] ^ DATA[43] ^ DATA[44] ^ DATA[46] ^ DATA[47] ^ DATA[51] ^ DATA[52] ^ DATA[53] ^ DATA[55] ^ DATA[58] ^ DATA[60] ^ DATA[61] ^ DATA[64] ^ DATA[66] ^ DATA[67] ^ DATA[68] ^ DATA[69] ^ DATA[70] ^ DATA[71] ^ DATA[74] ^ DATA[76] ^ DATA[77] ^ DATA[78] ^ DATA[79] ^ DATA[80] ^ DATA[81] ^ DATA[83] ^ DATA[84] ^ DATA[85] ^ DATA[86] ^ DATA[88] ^ DATA[89] ^ DATA[96] ^ DATA[98] ^ DATA[102] ^ DATA[104] ^ DATA[106] ^ DATA[108] ^ DATA[110] ^ DATA[113] ^ DATA[114] ^ DATA[115] ^ DATA[117] ^ DATA[119] ^ DATA[120] ^ DATA[121] ^ DATA[127] ^ DATA[129] ^ DATA[131] ^ DATA[136] ^ DATA[138] ^ DATA[140] ^ DATA[142] ^ DATA[143];
  assign CRC_OUT[10] = CRC_IN[1] ^ CRC_IN[3] ^ CRC_IN[5] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[18] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[27] ^ CRC_IN[29] ^ DATA[0] ^ DATA[2] ^ DATA[3] ^ DATA[5] ^ DATA[9] ^ DATA[13] ^ DATA[14] ^ DATA[16] ^ DATA[19] ^ DATA[26] ^ DATA[28] ^ DATA[29] ^ DATA[31] ^ DATA[32] ^ DATA[33] ^ DATA[35] ^ DATA[36] ^ DATA[39] ^ DATA[40] ^ DATA[42] ^ DATA[50] ^ DATA[52] ^ DATA[55] ^ DATA[56] ^ DATA[58] ^ DATA[59] ^ DATA[60] ^ DATA[62] ^ DATA[63] ^ DATA[66] ^ DATA[69] ^ DATA[70] ^ DATA[71] ^ DATA[73] ^ DATA[75] ^ DATA[77] ^ DATA[78] ^ DATA[80] ^ DATA[83] ^ DATA[86] ^ DATA[89] ^ DATA[90] ^ DATA[94] ^ DATA[95] ^ DATA[96] ^ DATA[98] ^ DATA[101] ^ DATA[104] ^ DATA[105] ^ DATA[106] ^ DATA[107] ^ DATA[109] ^ DATA[110] ^ DATA[113] ^ DATA[115] ^ DATA[117] ^ DATA[119] ^ DATA[120] ^ DATA[121] ^ DATA[122] ^ DATA[123] ^ DATA[125] ^ DATA[126] ^ DATA[127] ^ DATA[130] ^ DATA[134] ^ DATA[135] ^ DATA[136] ^ DATA[139] ^ DATA[141];
  assign CRC_OUT[11] = CRC_IN[1] ^ CRC_IN[5] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[22] ^ CRC_IN[28] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[0] ^ DATA[1] ^ DATA[3] ^ DATA[4] ^ DATA[9] ^ DATA[12] ^ DATA[14] ^ DATA[15] ^ DATA[16] ^ DATA[17] ^ DATA[20] ^ DATA[24] ^ DATA[25] ^ DATA[26] ^ DATA[27] ^ DATA[28] ^ DATA[31] ^ DATA[33] ^ DATA[36] ^ DATA[40] ^ DATA[41] ^ DATA[43] ^ DATA[44] ^ DATA[45] ^ DATA[47] ^ DATA[48] ^ DATA[50] ^ DATA[51] ^ DATA[54] ^ DATA[55] ^ DATA[56] ^ DATA[57] ^ DATA[58] ^ DATA[59] ^ DATA[64] ^ DATA[65] ^ DATA[66] ^ DATA[68] ^ DATA[70] ^ DATA[71] ^ DATA[73] ^ DATA[74] ^ DATA[76] ^ DATA[78] ^ DATA[82] ^ DATA[83] ^ DATA[85] ^ DATA[90] ^ DATA[91] ^ DATA[94] ^ DATA[98] ^ DATA[101] ^ DATA[102] ^ DATA[103] ^ DATA[104] ^ DATA[105] ^ DATA[107] ^ DATA[108] ^ DATA[113] ^ DATA[117] ^ DATA[119] ^ DATA[120] ^ DATA[121] ^ DATA[122] ^ DATA[124] ^ DATA[125] ^ DATA[131] ^ DATA[132] ^ DATA[134] ^ DATA[140] ^ DATA[142] ^ DATA[143];
  assign CRC_OUT[12] = CRC_IN[1] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[29] ^ DATA[0] ^ DATA[1] ^ DATA[2] ^ DATA[4] ^ DATA[5] ^ DATA[6] ^ DATA[9] ^ DATA[12] ^ DATA[13] ^ DATA[15] ^ DATA[17] ^ DATA[18] ^ DATA[21] ^ DATA[24] ^ DATA[27] ^ DATA[30] ^ DATA[31] ^ DATA[41] ^ DATA[42] ^ DATA[46] ^ DATA[47] ^ DATA[49] ^ DATA[50] ^ DATA[51] ^ DATA[52] ^ DATA[53] ^ DATA[54] ^ DATA[56] ^ DATA[57] ^ DATA[59] ^ DATA[61] ^ DATA[63] ^ DATA[68] ^ DATA[69] ^ DATA[71] ^ DATA[73] ^ DATA[74] ^ DATA[75] ^ DATA[77] ^ DATA[81] ^ DATA[82] ^ DATA[85] ^ DATA[86] ^ DATA[87] ^ DATA[91] ^ DATA[92] ^ DATA[94] ^ DATA[96] ^ DATA[97] ^ DATA[98] ^ DATA[101] ^ DATA[102] ^ DATA[105] ^ DATA[108] ^ DATA[109] ^ DATA[110] ^ DATA[111] ^ DATA[113] ^ DATA[116] ^ DATA[117] ^ DATA[119] ^ DATA[120] ^ DATA[121] ^ DATA[122] ^ DATA[127] ^ DATA[128] ^ DATA[133] ^ DATA[134] ^ DATA[136] ^ DATA[137] ^ DATA[141];
  assign CRC_OUT[13] = CRC_IN[0] ^ CRC_IN[2] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[30] ^ DATA[1] ^ DATA[2] ^ DATA[3] ^ DATA[5] ^ DATA[6] ^ DATA[7] ^ DATA[10] ^ DATA[13] ^ DATA[14] ^ DATA[16] ^ DATA[18] ^ DATA[19] ^ DATA[22] ^ DATA[25] ^ DATA[28] ^ DATA[31] ^ DATA[32] ^ DATA[42] ^ DATA[43] ^ DATA[47] ^ DATA[48] ^ DATA[50] ^ DATA[51] ^ DATA[52] ^ DATA[53] ^ DATA[54] ^ DATA[55] ^ DATA[57] ^ DATA[58] ^ DATA[60] ^ DATA[62] ^ DATA[64] ^ DATA[69] ^ DATA[70] ^ DATA[72] ^ DATA[74] ^ DATA[75] ^ DATA[76] ^ DATA[78] ^ DATA[82] ^ DATA[83] ^ DATA[86] ^ DATA[87] ^ DATA[88] ^ DATA[92] ^ DATA[93] ^ DATA[95] ^ DATA[97] ^ DATA[98] ^ DATA[99] ^ DATA[102] ^ DATA[103] ^ DATA[106] ^ DATA[109] ^ DATA[110] ^ DATA[111] ^ DATA[112] ^ DATA[114] ^ DATA[117] ^ DATA[118] ^ DATA[120] ^ DATA[121] ^ DATA[122] ^ DATA[123] ^ DATA[128] ^ DATA[129] ^ DATA[134] ^ DATA[135] ^ DATA[137] ^ DATA[138] ^ DATA[142];
  assign CRC_OUT[14] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[3] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[31] ^ DATA[2] ^ DATA[3] ^ DATA[4] ^ DATA[6] ^ DATA[7] ^ DATA[8] ^ DATA[11] ^ DATA[14] ^ DATA[15] ^ DATA[17] ^ DATA[19] ^ DATA[20] ^ DATA[23] ^ DATA[26] ^ DATA[29] ^ DATA[32] ^ DATA[33] ^ DATA[43] ^ DATA[44] ^ DATA[48] ^ DATA[49] ^ DATA[51] ^ DATA[52] ^ DATA[53] ^ DATA[54] ^ DATA[55] ^ DATA[56] ^ DATA[58] ^ DATA[59] ^ DATA[61] ^ DATA[63] ^ DATA[65] ^ DATA[70] ^ DATA[71] ^ DATA[73] ^ DATA[75] ^ DATA[76] ^ DATA[77] ^ DATA[79] ^ DATA[83] ^ DATA[84] ^ DATA[87] ^ DATA[88] ^ DATA[89] ^ DATA[93] ^ DATA[94] ^ DATA[96] ^ DATA[98] ^ DATA[99] ^ DATA[100] ^ DATA[103] ^ DATA[104] ^ DATA[107] ^ DATA[110] ^ DATA[111] ^ DATA[112] ^ DATA[113] ^ DATA[115] ^ DATA[118] ^ DATA[119] ^ DATA[121] ^ DATA[122] ^ DATA[123] ^ DATA[124] ^ DATA[129] ^ DATA[130] ^ DATA[135] ^ DATA[136] ^ DATA[138] ^ DATA[139] ^ DATA[143];
  assign CRC_OUT[15] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[4] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[27] ^ CRC_IN[28] ^ DATA[3] ^ DATA[4] ^ DATA[5] ^ DATA[7] ^ DATA[8] ^ DATA[9] ^ DATA[12] ^ DATA[15] ^ DATA[16] ^ DATA[18] ^ DATA[20] ^ DATA[21] ^ DATA[24] ^ DATA[27] ^ DATA[30] ^ DATA[33] ^ DATA[34] ^ DATA[44] ^ DATA[45] ^ DATA[49] ^ DATA[50] ^ DATA[52] ^ DATA[53] ^ DATA[54] ^ DATA[55] ^ DATA[56] ^ DATA[57] ^ DATA[59] ^ DATA[60] ^ DATA[62] ^ DATA[64] ^ DATA[66] ^ DATA[71] ^ DATA[72] ^ DATA[74] ^ DATA[76] ^ DATA[77] ^ DATA[78] ^ DATA[80] ^ DATA[84] ^ DATA[85] ^ DATA[88] ^ DATA[89] ^ DATA[90] ^ DATA[94] ^ DATA[95] ^ DATA[97] ^ DATA[99] ^ DATA[100] ^ DATA[101] ^ DATA[104] ^ DATA[105] ^ DATA[108] ^ DATA[111] ^ DATA[112] ^ DATA[113] ^ DATA[114] ^ DATA[116] ^ DATA[119] ^ DATA[120] ^ DATA[122] ^ DATA[123] ^ DATA[124] ^ DATA[125] ^ DATA[130] ^ DATA[131] ^ DATA[136] ^ DATA[137] ^ DATA[139] ^ DATA[140];
  assign CRC_OUT[16] = CRC_IN[0] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[12] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[19] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[26] ^ CRC_IN[28] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[0] ^ DATA[4] ^ DATA[5] ^ DATA[8] ^ DATA[12] ^ DATA[13] ^ DATA[17] ^ DATA[19] ^ DATA[21] ^ DATA[22] ^ DATA[24] ^ DATA[26] ^ DATA[29] ^ DATA[30] ^ DATA[32] ^ DATA[35] ^ DATA[37] ^ DATA[44] ^ DATA[46] ^ DATA[47] ^ DATA[48] ^ DATA[51] ^ DATA[56] ^ DATA[57] ^ DATA[66] ^ DATA[68] ^ DATA[75] ^ DATA[77] ^ DATA[78] ^ DATA[82] ^ DATA[83] ^ DATA[84] ^ DATA[86] ^ DATA[87] ^ DATA[89] ^ DATA[90] ^ DATA[91] ^ DATA[94] ^ DATA[97] ^ DATA[99] ^ DATA[100] ^ DATA[102] ^ DATA[103] ^ DATA[104] ^ DATA[105] ^ DATA[109] ^ DATA[110] ^ DATA[111] ^ DATA[112] ^ DATA[115] ^ DATA[116] ^ DATA[118] ^ DATA[119] ^ DATA[120] ^ DATA[121] ^ DATA[124] ^ DATA[127] ^ DATA[128] ^ DATA[131] ^ DATA[134] ^ DATA[135] ^ DATA[136] ^ DATA[138] ^ DATA[140] ^ DATA[141] ^ DATA[143];
  assign CRC_OUT[17] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[13] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[20] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[27] ^ CRC_IN[29] ^ CRC_IN[30] ^ DATA[1] ^ DATA[5] ^ DATA[6] ^ DATA[9] ^ DATA[13] ^ DATA[14] ^ DATA[18] ^ DATA[20] ^ DATA[22] ^ DATA[23] ^ DATA[25] ^ DATA[27] ^ DATA[30] ^ DATA[31] ^ DATA[33] ^ DATA[36] ^ DATA[38] ^ DATA[45] ^ DATA[47] ^ DATA[48] ^ DATA[49] ^ DATA[52] ^ DATA[57] ^ DATA[58] ^ DATA[67] ^ DATA[69] ^ DATA[76] ^ DATA[78] ^ DATA[79] ^ DATA[83] ^ DATA[84] ^ DATA[85] ^ DATA[87] ^ DATA[88] ^ DATA[90] ^ DATA[91] ^ DATA[92] ^ DATA[95] ^ DATA[98] ^ DATA[100] ^ DATA[101] ^ DATA[103] ^ DATA[104] ^ DATA[105] ^ DATA[106] ^ DATA[110] ^ DATA[111] ^ DATA[112] ^ DATA[113] ^ DATA[116] ^ DATA[117] ^ DATA[119] ^ DATA[120] ^ DATA[121] ^ DATA[122] ^ DATA[125] ^ DATA[128] ^ DATA[129] ^ DATA[132] ^ DATA[135] ^ DATA[136] ^ DATA[137] ^ DATA[139] ^ DATA[141] ^ DATA[142];
  assign CRC_OUT[18] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[14] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[21] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[28] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[2] ^ DATA[6] ^ DATA[7] ^ DATA[10] ^ DATA[14] ^ DATA[15] ^ DATA[19] ^ DATA[21] ^ DATA[23] ^ DATA[24] ^ DATA[26] ^ DATA[28] ^ DATA[31] ^ DATA[32] ^ DATA[34] ^ DATA[37] ^ DATA[39] ^ DATA[46] ^ DATA[48] ^ DATA[49] ^ DATA[50] ^ DATA[53] ^ DATA[58] ^ DATA[59] ^ DATA[68] ^ DATA[70] ^ DATA[77] ^ DATA[79] ^ DATA[80] ^ DATA[84] ^ DATA[85] ^ DATA[86] ^ DATA[88] ^ DATA[89] ^ DATA[91] ^ DATA[92] ^ DATA[93] ^ DATA[96] ^ DATA[99] ^ DATA[101] ^ DATA[102] ^ DATA[104] ^ DATA[105] ^ DATA[106] ^ DATA[107] ^ DATA[111] ^ DATA[112] ^ DATA[113] ^ DATA[114] ^ DATA[117] ^ DATA[118] ^ DATA[120] ^ DATA[121] ^ DATA[122] ^ DATA[123] ^ DATA[126] ^ DATA[129] ^ DATA[130] ^ DATA[133] ^ DATA[136] ^ DATA[137] ^ DATA[138] ^ DATA[140] ^ DATA[142] ^ DATA[143];
  assign CRC_OUT[19] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[15] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[22] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[3] ^ DATA[7] ^ DATA[8] ^ DATA[11] ^ DATA[15] ^ DATA[16] ^ DATA[20] ^ DATA[22] ^ DATA[24] ^ DATA[25] ^ DATA[27] ^ DATA[29] ^ DATA[32] ^ DATA[33] ^ DATA[35] ^ DATA[38] ^ DATA[40] ^ DATA[47] ^ DATA[49] ^ DATA[50] ^ DATA[51] ^ DATA[54] ^ DATA[59] ^ DATA[60] ^ DATA[69] ^ DATA[71] ^ DATA[78] ^ DATA[80] ^ DATA[81] ^ DATA[85] ^ DATA[86] ^ DATA[87] ^ DATA[89] ^ DATA[90] ^ DATA[92] ^ DATA[93] ^ DATA[94] ^ DATA[97] ^ DATA[100] ^ DATA[102] ^ DATA[103] ^ DATA[105] ^ DATA[106] ^ DATA[107] ^ DATA[108] ^ DATA[112] ^ DATA[113] ^ DATA[114] ^ DATA[115] ^ DATA[118] ^ DATA[119] ^ DATA[121] ^ DATA[122] ^ DATA[123] ^ DATA[124] ^ DATA[127] ^ DATA[130] ^ DATA[131] ^ DATA[134] ^ DATA[137] ^ DATA[138] ^ DATA[139] ^ DATA[141] ^ DATA[143];
  assign CRC_OUT[20] = CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[16] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[23] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[28] ^ CRC_IN[30] ^ DATA[4] ^ DATA[8] ^ DATA[9] ^ DATA[12] ^ DATA[16] ^ DATA[17] ^ DATA[21] ^ DATA[23] ^ DATA[25] ^ DATA[26] ^ DATA[28] ^ DATA[30] ^ DATA[33] ^ DATA[34] ^ DATA[36] ^ DATA[39] ^ DATA[41] ^ DATA[48] ^ DATA[50] ^ DATA[51] ^ DATA[52] ^ DATA[55] ^ DATA[60] ^ DATA[61] ^ DATA[70] ^ DATA[72] ^ DATA[79] ^ DATA[81] ^ DATA[82] ^ DATA[86] ^ DATA[87] ^ DATA[88] ^ DATA[90] ^ DATA[91] ^ DATA[93] ^ DATA[94] ^ DATA[95] ^ DATA[98] ^ DATA[101] ^ DATA[103] ^ DATA[104] ^ DATA[106] ^ DATA[107] ^ DATA[108] ^ DATA[109] ^ DATA[113] ^ DATA[114] ^ DATA[115] ^ DATA[116] ^ DATA[119] ^ DATA[120] ^ DATA[122] ^ DATA[123] ^ DATA[124] ^ DATA[125] ^ DATA[128] ^ DATA[131] ^ DATA[132] ^ DATA[135] ^ DATA[138] ^ DATA[139] ^ DATA[140] ^ DATA[142];
  assign CRC_OUT[21] = CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[17] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[24] ^ CRC_IN[27] ^ CRC_IN[28] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[5] ^ DATA[9] ^ DATA[10] ^ DATA[13] ^ DATA[17] ^ DATA[18] ^ DATA[22] ^ DATA[24] ^ DATA[26] ^ DATA[27] ^ DATA[29] ^ DATA[31] ^ DATA[34] ^ DATA[35] ^ DATA[37] ^ DATA[40] ^ DATA[42] ^ DATA[49] ^ DATA[51] ^ DATA[52] ^ DATA[53] ^ DATA[56] ^ DATA[61] ^ DATA[62] ^ DATA[71] ^ DATA[73] ^ DATA[80] ^ DATA[82] ^ DATA[83] ^ DATA[87] ^ DATA[88] ^ DATA[89] ^ DATA[91] ^ DATA[92] ^ DATA[94] ^ DATA[95] ^ DATA[96] ^ DATA[99] ^ DATA[102] ^ DATA[104] ^ DATA[105] ^ DATA[107] ^ DATA[108] ^ DATA[109] ^ DATA[110] ^ DATA[114] ^ DATA[115] ^ DATA[116] ^ DATA[117] ^ DATA[120] ^ DATA[121] ^ DATA[123] ^ DATA[124] ^ DATA[125] ^ DATA[126] ^ DATA[129] ^ DATA[132] ^ DATA[133] ^ DATA[136] ^ DATA[139] ^ DATA[140] ^ DATA[141] ^ DATA[143];
  assign CRC_OUT[22] = CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[7] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[16] ^ CRC_IN[18] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[28] ^ CRC_IN[29] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[0] ^ DATA[9] ^ DATA[11] ^ DATA[12] ^ DATA[14] ^ DATA[16] ^ DATA[18] ^ DATA[19] ^ DATA[23] ^ DATA[24] ^ DATA[26] ^ DATA[27] ^ DATA[29] ^ DATA[31] ^ DATA[34] ^ DATA[35] ^ DATA[36] ^ DATA[37] ^ DATA[38] ^ DATA[41] ^ DATA[43] ^ DATA[44] ^ DATA[45] ^ DATA[47] ^ DATA[48] ^ DATA[52] ^ DATA[55] ^ DATA[57] ^ DATA[58] ^ DATA[60] ^ DATA[61] ^ DATA[62] ^ DATA[65] ^ DATA[66] ^ DATA[67] ^ DATA[68] ^ DATA[73] ^ DATA[74] ^ DATA[79] ^ DATA[82] ^ DATA[85] ^ DATA[87] ^ DATA[88] ^ DATA[89] ^ DATA[90] ^ DATA[92] ^ DATA[93] ^ DATA[94] ^ DATA[98] ^ DATA[99] ^ DATA[100] ^ DATA[101] ^ DATA[104] ^ DATA[105] ^ DATA[108] ^ DATA[109] ^ DATA[113] ^ DATA[114] ^ DATA[115] ^ DATA[119] ^ DATA[121] ^ DATA[122] ^ DATA[123] ^ DATA[124] ^ DATA[128] ^ DATA[130] ^ DATA[132] ^ DATA[133] ^ DATA[135] ^ DATA[136] ^ DATA[140] ^ DATA[141] ^ DATA[142] ^ DATA[143];
  assign CRC_OUT[23] = CRC_IN[1] ^ CRC_IN[3] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[23] ^ CRC_IN[29] ^ CRC_IN[30] ^ DATA[0] ^ DATA[1] ^ DATA[6] ^ DATA[9] ^ DATA[13] ^ DATA[15] ^ DATA[16] ^ DATA[17] ^ DATA[19] ^ DATA[20] ^ DATA[26] ^ DATA[27] ^ DATA[29] ^ DATA[31] ^ DATA[34] ^ DATA[35] ^ DATA[36] ^ DATA[38] ^ DATA[39] ^ DATA[42] ^ DATA[46] ^ DATA[47] ^ DATA[49] ^ DATA[50] ^ DATA[54] ^ DATA[55] ^ DATA[56] ^ DATA[59] ^ DATA[60] ^ DATA[62] ^ DATA[65] ^ DATA[69] ^ DATA[72] ^ DATA[73] ^ DATA[74] ^ DATA[75] ^ DATA[79] ^ DATA[80] ^ DATA[81] ^ DATA[82] ^ DATA[84] ^ DATA[85] ^ DATA[86] ^ DATA[87] ^ DATA[88] ^ DATA[89] ^ DATA[90] ^ DATA[91] ^ DATA[93] ^ DATA[96] ^ DATA[97] ^ DATA[98] ^ DATA[100] ^ DATA[102] ^ DATA[103] ^ DATA[104] ^ DATA[105] ^ DATA[109] ^ DATA[111] ^ DATA[113] ^ DATA[115] ^ DATA[117] ^ DATA[118] ^ DATA[119] ^ DATA[120] ^ DATA[122] ^ DATA[124] ^ DATA[126] ^ DATA[127] ^ DATA[128] ^ DATA[129] ^ DATA[131] ^ DATA[132] ^ DATA[133] ^ DATA[135] ^ DATA[141] ^ DATA[142];
  assign CRC_OUT[24] = CRC_IN[0] ^ CRC_IN[2] ^ CRC_IN[4] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[11] ^ CRC_IN[13] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[24] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[1] ^ DATA[2] ^ DATA[7] ^ DATA[10] ^ DATA[14] ^ DATA[16] ^ DATA[17] ^ DATA[18] ^ DATA[20] ^ DATA[21] ^ DATA[27] ^ DATA[28] ^ DATA[30] ^ DATA[32] ^ DATA[35] ^ DATA[36] ^ DATA[37] ^ DATA[39] ^ DATA[40] ^ DATA[43] ^ DATA[47] ^ DATA[48] ^ DATA[50] ^ DATA[51] ^ DATA[55] ^ DATA[56] ^ DATA[57] ^ DATA[60] ^ DATA[61] ^ DATA[63] ^ DATA[66] ^ DATA[70] ^ DATA[73] ^ DATA[74] ^ DATA[75] ^ DATA[76] ^ DATA[80] ^ DATA[81] ^ DATA[82] ^ DATA[83] ^ DATA[85] ^ DATA[86] ^ DATA[87] ^ DATA[88] ^ DATA[89] ^ DATA[90] ^ DATA[91] ^ DATA[92] ^ DATA[94] ^ DATA[97] ^ DATA[98] ^ DATA[99] ^ DATA[101] ^ DATA[103] ^ DATA[104] ^ DATA[105] ^ DATA[106] ^ DATA[110] ^ DATA[112] ^ DATA[114] ^ DATA[116] ^ DATA[118] ^ DATA[119] ^ DATA[120] ^ DATA[121] ^ DATA[123] ^ DATA[125] ^ DATA[127] ^ DATA[128] ^ DATA[129] ^ DATA[130] ^ DATA[132] ^ DATA[133] ^ DATA[134] ^ DATA[136] ^ DATA[142] ^ DATA[143];
  assign CRC_OUT[25] = CRC_IN[1] ^ CRC_IN[3] ^ CRC_IN[5] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[14] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[25] ^ CRC_IN[31] ^ DATA[2] ^ DATA[3] ^ DATA[8] ^ DATA[11] ^ DATA[15] ^ DATA[17] ^ DATA[18] ^ DATA[19] ^ DATA[21] ^ DATA[22] ^ DATA[28] ^ DATA[29] ^ DATA[31] ^ DATA[33] ^ DATA[36] ^ DATA[37] ^ DATA[38] ^ DATA[40] ^ DATA[41] ^ DATA[44] ^ DATA[48] ^ DATA[49] ^ DATA[51] ^ DATA[52] ^ DATA[56] ^ DATA[57] ^ DATA[58] ^ DATA[61] ^ DATA[62] ^ DATA[64] ^ DATA[67] ^ DATA[71] ^ DATA[74] ^ DATA[75] ^ DATA[76] ^ DATA[77] ^ DATA[81] ^ DATA[82] ^ DATA[83] ^ DATA[84] ^ DATA[86] ^ DATA[87] ^ DATA[88] ^ DATA[89] ^ DATA[90] ^ DATA[91] ^ DATA[92] ^ DATA[93] ^ DATA[95] ^ DATA[98] ^ DATA[99] ^ DATA[100] ^ DATA[102] ^ DATA[104] ^ DATA[105] ^ DATA[106] ^ DATA[107] ^ DATA[111] ^ DATA[113] ^ DATA[115] ^ DATA[117] ^ DATA[119] ^ DATA[120] ^ DATA[121] ^ DATA[122] ^ DATA[124] ^ DATA[126] ^ DATA[128] ^ DATA[129] ^ DATA[130] ^ DATA[131] ^ DATA[133] ^ DATA[134] ^ DATA[135] ^ DATA[137] ^ DATA[143];
  assign CRC_OUT[26] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[5] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[14] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[31] ^ DATA[0] ^ DATA[3] ^ DATA[4] ^ DATA[6] ^ DATA[10] ^ DATA[18] ^ DATA[19] ^ DATA[20] ^ DATA[22] ^ DATA[23] ^ DATA[24] ^ DATA[25] ^ DATA[26] ^ DATA[28] ^ DATA[31] ^ DATA[38] ^ DATA[39] ^ DATA[41] ^ DATA[42] ^ DATA[44] ^ DATA[47] ^ DATA[48] ^ DATA[49] ^ DATA[52] ^ DATA[54] ^ DATA[55] ^ DATA[57] ^ DATA[59] ^ DATA[60] ^ DATA[61] ^ DATA[62] ^ DATA[66] ^ DATA[67] ^ DATA[73] ^ DATA[75] ^ DATA[76] ^ DATA[77] ^ DATA[78] ^ DATA[79] ^ DATA[81] ^ DATA[88] ^ DATA[89] ^ DATA[90] ^ DATA[91] ^ DATA[92] ^ DATA[93] ^ DATA[95] ^ DATA[97] ^ DATA[98] ^ DATA[100] ^ DATA[104] ^ DATA[105] ^ DATA[107] ^ DATA[108] ^ DATA[110] ^ DATA[111] ^ DATA[112] ^ DATA[113] ^ DATA[117] ^ DATA[119] ^ DATA[120] ^ DATA[121] ^ DATA[122] ^ DATA[126] ^ DATA[128] ^ DATA[129] ^ DATA[130] ^ DATA[131] ^ DATA[137] ^ DATA[138] ^ DATA[143];
  assign CRC_OUT[27] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[6] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[15] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[26] ^ CRC_IN[27] ^ DATA[1] ^ DATA[4] ^ DATA[5] ^ DATA[7] ^ DATA[11] ^ DATA[19] ^ DATA[20] ^ DATA[21] ^ DATA[23] ^ DATA[24] ^ DATA[25] ^ DATA[26] ^ DATA[27] ^ DATA[29] ^ DATA[32] ^ DATA[39] ^ DATA[40] ^ DATA[42] ^ DATA[43] ^ DATA[45] ^ DATA[48] ^ DATA[49] ^ DATA[50] ^ DATA[53] ^ DATA[55] ^ DATA[56] ^ DATA[58] ^ DATA[60] ^ DATA[61] ^ DATA[62] ^ DATA[63] ^ DATA[67] ^ DATA[68] ^ DATA[74] ^ DATA[76] ^ DATA[77] ^ DATA[78] ^ DATA[79] ^ DATA[80] ^ DATA[82] ^ DATA[89] ^ DATA[90] ^ DATA[91] ^ DATA[92] ^ DATA[93] ^ DATA[94] ^ DATA[96] ^ DATA[98] ^ DATA[99] ^ DATA[101] ^ DATA[105] ^ DATA[106] ^ DATA[108] ^ DATA[109] ^ DATA[111] ^ DATA[112] ^ DATA[113] ^ DATA[114] ^ DATA[118] ^ DATA[120] ^ DATA[121] ^ DATA[122] ^ DATA[123] ^ DATA[127] ^ DATA[129] ^ DATA[130] ^ DATA[131] ^ DATA[132] ^ DATA[138] ^ DATA[139];
  assign CRC_OUT[28] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[7] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[16] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[27] ^ CRC_IN[28] ^ DATA[2] ^ DATA[5] ^ DATA[6] ^ DATA[8] ^ DATA[12] ^ DATA[20] ^ DATA[21] ^ DATA[22] ^ DATA[24] ^ DATA[25] ^ DATA[26] ^ DATA[27] ^ DATA[28] ^ DATA[30] ^ DATA[33] ^ DATA[40] ^ DATA[41] ^ DATA[43] ^ DATA[44] ^ DATA[46] ^ DATA[49] ^ DATA[50] ^ DATA[51] ^ DATA[54] ^ DATA[56] ^ DATA[57] ^ DATA[59] ^ DATA[61] ^ DATA[62] ^ DATA[63] ^ DATA[64] ^ DATA[68] ^ DATA[69] ^ DATA[75] ^ DATA[77] ^ DATA[78] ^ DATA[79] ^ DATA[80] ^ DATA[81] ^ DATA[83] ^ DATA[90] ^ DATA[91] ^ DATA[92] ^ DATA[93] ^ DATA[94] ^ DATA[95] ^ DATA[97] ^ DATA[99] ^ DATA[100] ^ DATA[102] ^ DATA[106] ^ DATA[107] ^ DATA[109] ^ DATA[110] ^ DATA[112] ^ DATA[113] ^ DATA[114] ^ DATA[115] ^ DATA[119] ^ DATA[121] ^ DATA[122] ^ DATA[123] ^ DATA[124] ^ DATA[128] ^ DATA[130] ^ DATA[131] ^ DATA[132] ^ DATA[133] ^ DATA[139] ^ DATA[140];
  assign CRC_OUT[29] = CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[17] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[28] ^ CRC_IN[29] ^ DATA[3] ^ DATA[6] ^ DATA[7] ^ DATA[9] ^ DATA[13] ^ DATA[21] ^ DATA[22] ^ DATA[23] ^ DATA[25] ^ DATA[26] ^ DATA[27] ^ DATA[28] ^ DATA[29] ^ DATA[31] ^ DATA[34] ^ DATA[41] ^ DATA[42] ^ DATA[44] ^ DATA[45] ^ DATA[47] ^ DATA[50] ^ DATA[51] ^ DATA[52] ^ DATA[55] ^ DATA[57] ^ DATA[58] ^ DATA[60] ^ DATA[62] ^ DATA[63] ^ DATA[64] ^ DATA[65] ^ DATA[69] ^ DATA[70] ^ DATA[76] ^ DATA[78] ^ DATA[79] ^ DATA[80] ^ DATA[81] ^ DATA[82] ^ DATA[84] ^ DATA[91] ^ DATA[92] ^ DATA[93] ^ DATA[94] ^ DATA[95] ^ DATA[96] ^ DATA[98] ^ DATA[100] ^ DATA[101] ^ DATA[103] ^ DATA[107] ^ DATA[108] ^ DATA[110] ^ DATA[111] ^ DATA[113] ^ DATA[114] ^ DATA[115] ^ DATA[116] ^ DATA[120] ^ DATA[122] ^ DATA[123] ^ DATA[124] ^ DATA[125] ^ DATA[129] ^ DATA[131] ^ DATA[132] ^ DATA[133] ^ DATA[134] ^ DATA[140] ^ DATA[141];
  assign CRC_OUT[30] = CRC_IN[0] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[9] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[18] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[29] ^ CRC_IN[30] ^ DATA[4] ^ DATA[7] ^ DATA[8] ^ DATA[10] ^ DATA[14] ^ DATA[22] ^ DATA[23] ^ DATA[24] ^ DATA[26] ^ DATA[27] ^ DATA[28] ^ DATA[29] ^ DATA[30] ^ DATA[32] ^ DATA[35] ^ DATA[42] ^ DATA[43] ^ DATA[45] ^ DATA[46] ^ DATA[48] ^ DATA[51] ^ DATA[52] ^ DATA[53] ^ DATA[56] ^ DATA[58] ^ DATA[59] ^ DATA[61] ^ DATA[63] ^ DATA[64] ^ DATA[65] ^ DATA[66] ^ DATA[70] ^ DATA[71] ^ DATA[77] ^ DATA[79] ^ DATA[80] ^ DATA[81] ^ DATA[82] ^ DATA[83] ^ DATA[85] ^ DATA[92] ^ DATA[93] ^ DATA[94] ^ DATA[95] ^ DATA[96] ^ DATA[97] ^ DATA[99] ^ DATA[101] ^ DATA[102] ^ DATA[104] ^ DATA[108] ^ DATA[109] ^ DATA[111] ^ DATA[112] ^ DATA[114] ^ DATA[115] ^ DATA[116] ^ DATA[117] ^ DATA[121] ^ DATA[123] ^ DATA[124] ^ DATA[125] ^ DATA[126] ^ DATA[130] ^ DATA[132] ^ DATA[133] ^ DATA[134] ^ DATA[135] ^ DATA[141] ^ DATA[142];
  assign CRC_OUT[31] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[19] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[5] ^ DATA[8] ^ DATA[9] ^ DATA[11] ^ DATA[15] ^ DATA[23] ^ DATA[24] ^ DATA[25] ^ DATA[27] ^ DATA[28] ^ DATA[29] ^ DATA[30] ^ DATA[31] ^ DATA[33] ^ DATA[36] ^ DATA[43] ^ DATA[44] ^ DATA[46] ^ DATA[47] ^ DATA[49] ^ DATA[52] ^ DATA[53] ^ DATA[54] ^ DATA[57] ^ DATA[59] ^ DATA[60] ^ DATA[62] ^ DATA[64] ^ DATA[65] ^ DATA[66] ^ DATA[67] ^ DATA[71] ^ DATA[72] ^ DATA[78] ^ DATA[80] ^ DATA[81] ^ DATA[82] ^ DATA[83] ^ DATA[84] ^ DATA[86] ^ DATA[93] ^ DATA[94] ^ DATA[95] ^ DATA[96] ^ DATA[97] ^ DATA[98] ^ DATA[100] ^ DATA[102] ^ DATA[103] ^ DATA[105] ^ DATA[109] ^ DATA[110] ^ DATA[112] ^ DATA[113] ^ DATA[115] ^ DATA[116] ^ DATA[117] ^ DATA[118] ^ DATA[122] ^ DATA[124] ^ DATA[125] ^ DATA[126] ^ DATA[127] ^ DATA[131] ^ DATA[133] ^ DATA[134] ^ DATA[135] ^ DATA[136] ^ DATA[142] ^ DATA[143];
endmodule
