// CRC polynomial coefficients: x^32 + x^26 + x^23 + x^22 + x^16 + x^12 + x^11 + x^10 + x^8 + x^7 + x^5 + x^4 + x^2 + x + 1
//                              0x4C11DB7 (hex)
// CRC width:                   32 bits
// CRC shift direction:         left (big endian)
// Input word width:            48 bits
`default_nettype none
module CRC_32 (
    input  wire [31:0] CRC_IN,
    input  wire [47:0] DATA,
    output wire [31:0] CRC_OUT
);
  assign CRC_OUT[0] = CRC_IN[0] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[18] ^ CRC_IN[21] ^ CRC_IN[28] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[0] ^ DATA[6] ^ DATA[9] ^ DATA[10] ^ DATA[12] ^ DATA[16] ^ DATA[24] ^ DATA[25] ^ DATA[26] ^ DATA[28] ^ DATA[29] ^ DATA[30] ^ DATA[31] ^ DATA[32] ^ DATA[34] ^ DATA[37] ^ DATA[44] ^ DATA[45] ^ DATA[47];
  assign CRC_OUT[1] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[8] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[28] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[0] ^ DATA[1] ^ DATA[6] ^ DATA[7] ^ DATA[9] ^ DATA[11] ^ DATA[12] ^ DATA[13] ^ DATA[16] ^ DATA[17] ^ DATA[24] ^ DATA[27] ^ DATA[28] ^ DATA[33] ^ DATA[34] ^ DATA[35] ^ DATA[37] ^ DATA[38] ^ DATA[44] ^ DATA[46] ^ DATA[47];
  assign CRC_OUT[2] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[28] ^ DATA[0] ^ DATA[1] ^ DATA[2] ^ DATA[6] ^ DATA[7] ^ DATA[8] ^ DATA[9] ^ DATA[13] ^ DATA[14] ^ DATA[16] ^ DATA[17] ^ DATA[18] ^ DATA[24] ^ DATA[26] ^ DATA[30] ^ DATA[31] ^ DATA[32] ^ DATA[35] ^ DATA[36] ^ DATA[37] ^ DATA[38] ^ DATA[39] ^ DATA[44];
  assign CRC_OUT[3] = CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[9] ^ CRC_IN[11] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[29] ^ DATA[1] ^ DATA[2] ^ DATA[3] ^ DATA[7] ^ DATA[8] ^ DATA[9] ^ DATA[10] ^ DATA[14] ^ DATA[15] ^ DATA[17] ^ DATA[18] ^ DATA[19] ^ DATA[25] ^ DATA[27] ^ DATA[31] ^ DATA[32] ^ DATA[33] ^ DATA[36] ^ DATA[37] ^ DATA[38] ^ DATA[39] ^ DATA[40] ^ DATA[45];
  assign CRC_OUT[4] = CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[17] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[28] ^ CRC_IN[29] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[0] ^ DATA[2] ^ DATA[3] ^ DATA[4] ^ DATA[6] ^ DATA[8] ^ DATA[11] ^ DATA[12] ^ DATA[15] ^ DATA[18] ^ DATA[19] ^ DATA[20] ^ DATA[24] ^ DATA[25] ^ DATA[29] ^ DATA[30] ^ DATA[31] ^ DATA[33] ^ DATA[38] ^ DATA[39] ^ DATA[40] ^ DATA[41] ^ DATA[44] ^ DATA[45] ^ DATA[46] ^ DATA[47];
  assign CRC_OUT[5] = CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[8] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[21] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[28] ^ CRC_IN[30] ^ DATA[0] ^ DATA[1] ^ DATA[3] ^ DATA[4] ^ DATA[5] ^ DATA[6] ^ DATA[7] ^ DATA[10] ^ DATA[13] ^ DATA[19] ^ DATA[20] ^ DATA[21] ^ DATA[24] ^ DATA[28] ^ DATA[29] ^ DATA[37] ^ DATA[39] ^ DATA[40] ^ DATA[41] ^ DATA[42] ^ DATA[44] ^ DATA[46];
  assign CRC_OUT[6] = CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[9] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[22] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[1] ^ DATA[2] ^ DATA[4] ^ DATA[5] ^ DATA[6] ^ DATA[7] ^ DATA[8] ^ DATA[11] ^ DATA[14] ^ DATA[20] ^ DATA[21] ^ DATA[22] ^ DATA[25] ^ DATA[29] ^ DATA[30] ^ DATA[38] ^ DATA[40] ^ DATA[41] ^ DATA[42] ^ DATA[43] ^ DATA[45] ^ DATA[47];
  assign CRC_OUT[7] = CRC_IN[0] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[16] ^ CRC_IN[18] ^ CRC_IN[21] ^ CRC_IN[23] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[29] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[0] ^ DATA[2] ^ DATA[3] ^ DATA[5] ^ DATA[7] ^ DATA[8] ^ DATA[10] ^ DATA[15] ^ DATA[16] ^ DATA[21] ^ DATA[22] ^ DATA[23] ^ DATA[24] ^ DATA[25] ^ DATA[28] ^ DATA[29] ^ DATA[32] ^ DATA[34] ^ DATA[37] ^ DATA[39] ^ DATA[41] ^ DATA[42] ^ DATA[43] ^ DATA[45] ^ DATA[46] ^ DATA[47];
  assign CRC_OUT[8] = CRC_IN[1] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[12] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[24] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[29] ^ CRC_IN[30] ^ DATA[0] ^ DATA[1] ^ DATA[3] ^ DATA[4] ^ DATA[8] ^ DATA[10] ^ DATA[11] ^ DATA[12] ^ DATA[17] ^ DATA[22] ^ DATA[23] ^ DATA[28] ^ DATA[31] ^ DATA[32] ^ DATA[33] ^ DATA[34] ^ DATA[35] ^ DATA[37] ^ DATA[38] ^ DATA[40] ^ DATA[42] ^ DATA[43] ^ DATA[45] ^ DATA[46];
  assign CRC_OUT[9] = CRC_IN[2] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[13] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[25] ^ CRC_IN[27] ^ CRC_IN[28] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[1] ^ DATA[2] ^ DATA[4] ^ DATA[5] ^ DATA[9] ^ DATA[11] ^ DATA[12] ^ DATA[13] ^ DATA[18] ^ DATA[23] ^ DATA[24] ^ DATA[29] ^ DATA[32] ^ DATA[33] ^ DATA[34] ^ DATA[35] ^ DATA[36] ^ DATA[38] ^ DATA[39] ^ DATA[41] ^ DATA[43] ^ DATA[44] ^ DATA[46] ^ DATA[47];
  assign CRC_OUT[10] = CRC_IN[0] ^ CRC_IN[3] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[26] ^ DATA[0] ^ DATA[2] ^ DATA[3] ^ DATA[5] ^ DATA[9] ^ DATA[13] ^ DATA[14] ^ DATA[16] ^ DATA[19] ^ DATA[26] ^ DATA[28] ^ DATA[29] ^ DATA[31] ^ DATA[32] ^ DATA[33] ^ DATA[35] ^ DATA[36] ^ DATA[39] ^ DATA[40] ^ DATA[42];
  assign CRC_OUT[11] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[4] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[15] ^ CRC_IN[17] ^ CRC_IN[20] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[27] ^ CRC_IN[28] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[0] ^ DATA[1] ^ DATA[3] ^ DATA[4] ^ DATA[9] ^ DATA[12] ^ DATA[14] ^ DATA[15] ^ DATA[16] ^ DATA[17] ^ DATA[20] ^ DATA[24] ^ DATA[25] ^ DATA[26] ^ DATA[27] ^ DATA[28] ^ DATA[31] ^ DATA[33] ^ DATA[36] ^ DATA[40] ^ DATA[41] ^ DATA[43] ^ DATA[44] ^ DATA[45] ^ DATA[47];
  assign CRC_OUT[12] = CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[5] ^ CRC_IN[8] ^ CRC_IN[11] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[0] ^ DATA[1] ^ DATA[2] ^ DATA[4] ^ DATA[5] ^ DATA[6] ^ DATA[9] ^ DATA[12] ^ DATA[13] ^ DATA[15] ^ DATA[17] ^ DATA[18] ^ DATA[21] ^ DATA[24] ^ DATA[27] ^ DATA[30] ^ DATA[31] ^ DATA[41] ^ DATA[42] ^ DATA[46] ^ DATA[47];
  assign CRC_OUT[13] = CRC_IN[0] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[6] ^ CRC_IN[9] ^ CRC_IN[12] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[31] ^ DATA[1] ^ DATA[2] ^ DATA[3] ^ DATA[5] ^ DATA[6] ^ DATA[7] ^ DATA[10] ^ DATA[13] ^ DATA[14] ^ DATA[16] ^ DATA[18] ^ DATA[19] ^ DATA[22] ^ DATA[25] ^ DATA[28] ^ DATA[31] ^ DATA[32] ^ DATA[42] ^ DATA[43] ^ DATA[47];
  assign CRC_OUT[14] = CRC_IN[1] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[7] ^ CRC_IN[10] ^ CRC_IN[13] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[27] ^ CRC_IN[28] ^ DATA[2] ^ DATA[3] ^ DATA[4] ^ DATA[6] ^ DATA[7] ^ DATA[8] ^ DATA[11] ^ DATA[14] ^ DATA[15] ^ DATA[17] ^ DATA[19] ^ DATA[20] ^ DATA[23] ^ DATA[26] ^ DATA[29] ^ DATA[32] ^ DATA[33] ^ DATA[43] ^ DATA[44];
  assign CRC_OUT[15] = CRC_IN[0] ^ CRC_IN[2] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[8] ^ CRC_IN[11] ^ CRC_IN[14] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[28] ^ CRC_IN[29] ^ DATA[3] ^ DATA[4] ^ DATA[5] ^ DATA[7] ^ DATA[8] ^ DATA[9] ^ DATA[12] ^ DATA[15] ^ DATA[16] ^ DATA[18] ^ DATA[20] ^ DATA[21] ^ DATA[24] ^ DATA[27] ^ DATA[30] ^ DATA[33] ^ DATA[34] ^ DATA[44] ^ DATA[45];
  assign CRC_OUT[16] = CRC_IN[1] ^ CRC_IN[3] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[16] ^ CRC_IN[19] ^ CRC_IN[21] ^ CRC_IN[28] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[0] ^ DATA[4] ^ DATA[5] ^ DATA[8] ^ DATA[12] ^ DATA[13] ^ DATA[17] ^ DATA[19] ^ DATA[21] ^ DATA[22] ^ DATA[24] ^ DATA[26] ^ DATA[29] ^ DATA[30] ^ DATA[32] ^ DATA[35] ^ DATA[37] ^ DATA[44] ^ DATA[46] ^ DATA[47];
  assign CRC_OUT[17] = CRC_IN[2] ^ CRC_IN[4] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[9] ^ CRC_IN[11] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[17] ^ CRC_IN[20] ^ CRC_IN[22] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[1] ^ DATA[5] ^ DATA[6] ^ DATA[9] ^ DATA[13] ^ DATA[14] ^ DATA[18] ^ DATA[20] ^ DATA[22] ^ DATA[23] ^ DATA[25] ^ DATA[27] ^ DATA[30] ^ DATA[31] ^ DATA[33] ^ DATA[36] ^ DATA[38] ^ DATA[45] ^ DATA[47];
  assign CRC_OUT[18] = CRC_IN[3] ^ CRC_IN[5] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[15] ^ CRC_IN[16] ^ CRC_IN[18] ^ CRC_IN[21] ^ CRC_IN[23] ^ CRC_IN[30] ^ DATA[2] ^ DATA[6] ^ DATA[7] ^ DATA[10] ^ DATA[14] ^ DATA[15] ^ DATA[19] ^ DATA[21] ^ DATA[23] ^ DATA[24] ^ DATA[26] ^ DATA[28] ^ DATA[31] ^ DATA[32] ^ DATA[34] ^ DATA[37] ^ DATA[39] ^ DATA[46];
  assign CRC_OUT[19] = CRC_IN[0] ^ CRC_IN[4] ^ CRC_IN[6] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[11] ^ CRC_IN[13] ^ CRC_IN[16] ^ CRC_IN[17] ^ CRC_IN[19] ^ CRC_IN[22] ^ CRC_IN[24] ^ CRC_IN[31] ^ DATA[3] ^ DATA[7] ^ DATA[8] ^ DATA[11] ^ DATA[15] ^ DATA[16] ^ DATA[20] ^ DATA[22] ^ DATA[24] ^ DATA[25] ^ DATA[27] ^ DATA[29] ^ DATA[32] ^ DATA[33] ^ DATA[35] ^ DATA[38] ^ DATA[40] ^ DATA[47];
  assign CRC_OUT[20] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[5] ^ CRC_IN[7] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[14] ^ CRC_IN[17] ^ CRC_IN[18] ^ CRC_IN[20] ^ CRC_IN[23] ^ CRC_IN[25] ^ DATA[4] ^ DATA[8] ^ DATA[9] ^ DATA[12] ^ DATA[16] ^ DATA[17] ^ DATA[21] ^ DATA[23] ^ DATA[25] ^ DATA[26] ^ DATA[28] ^ DATA[30] ^ DATA[33] ^ DATA[34] ^ DATA[36] ^ DATA[39] ^ DATA[41];
  assign CRC_OUT[21] = CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[6] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[13] ^ CRC_IN[15] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[21] ^ CRC_IN[24] ^ CRC_IN[26] ^ DATA[5] ^ DATA[9] ^ DATA[10] ^ DATA[13] ^ DATA[17] ^ DATA[18] ^ DATA[22] ^ DATA[24] ^ DATA[26] ^ DATA[27] ^ DATA[29] ^ DATA[31] ^ DATA[34] ^ DATA[35] ^ DATA[37] ^ DATA[40] ^ DATA[42];
  assign CRC_OUT[22] = CRC_IN[0] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[13] ^ CRC_IN[15] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[25] ^ CRC_IN[27] ^ CRC_IN[28] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[0] ^ DATA[9] ^ DATA[11] ^ DATA[12] ^ DATA[14] ^ DATA[16] ^ DATA[18] ^ DATA[19] ^ DATA[23] ^ DATA[24] ^ DATA[26] ^ DATA[27] ^ DATA[29] ^ DATA[31] ^ DATA[34] ^ DATA[35] ^ DATA[36] ^ DATA[37] ^ DATA[38] ^ DATA[41] ^ DATA[43] ^ DATA[44] ^ DATA[45] ^ DATA[47];
  assign CRC_OUT[23] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[13] ^ CRC_IN[15] ^ CRC_IN[18] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[26] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[0] ^ DATA[1] ^ DATA[6] ^ DATA[9] ^ DATA[13] ^ DATA[15] ^ DATA[16] ^ DATA[17] ^ DATA[19] ^ DATA[20] ^ DATA[26] ^ DATA[27] ^ DATA[29] ^ DATA[31] ^ DATA[34] ^ DATA[35] ^ DATA[36] ^ DATA[38] ^ DATA[39] ^ DATA[42] ^ DATA[46] ^ DATA[47];
  assign CRC_OUT[24] = CRC_IN[0] ^ CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[14] ^ CRC_IN[16] ^ CRC_IN[19] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[27] ^ CRC_IN[31] ^ DATA[1] ^ DATA[2] ^ DATA[7] ^ DATA[10] ^ DATA[14] ^ DATA[16] ^ DATA[17] ^ DATA[18] ^ DATA[20] ^ DATA[21] ^ DATA[27] ^ DATA[28] ^ DATA[30] ^ DATA[32] ^ DATA[35] ^ DATA[36] ^ DATA[37] ^ DATA[39] ^ DATA[40] ^ DATA[43] ^ DATA[47];
  assign CRC_OUT[25] = CRC_IN[1] ^ CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[15] ^ CRC_IN[17] ^ CRC_IN[20] ^ CRC_IN[21] ^ CRC_IN[22] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[28] ^ DATA[2] ^ DATA[3] ^ DATA[8] ^ DATA[11] ^ DATA[15] ^ DATA[17] ^ DATA[18] ^ DATA[19] ^ DATA[21] ^ DATA[22] ^ DATA[28] ^ DATA[29] ^ DATA[31] ^ DATA[33] ^ DATA[36] ^ DATA[37] ^ DATA[38] ^ DATA[40] ^ DATA[41] ^ DATA[44];
  assign CRC_OUT[26] = CRC_IN[2] ^ CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[12] ^ CRC_IN[15] ^ CRC_IN[22] ^ CRC_IN[23] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[28] ^ CRC_IN[31] ^ DATA[0] ^ DATA[3] ^ DATA[4] ^ DATA[6] ^ DATA[10] ^ DATA[18] ^ DATA[19] ^ DATA[20] ^ DATA[22] ^ DATA[23] ^ DATA[24] ^ DATA[25] ^ DATA[26] ^ DATA[28] ^ DATA[31] ^ DATA[38] ^ DATA[39] ^ DATA[41] ^ DATA[42] ^ DATA[44] ^ DATA[47];
  assign CRC_OUT[27] = CRC_IN[3] ^ CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[13] ^ CRC_IN[16] ^ CRC_IN[23] ^ CRC_IN[24] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[29] ^ DATA[1] ^ DATA[4] ^ DATA[5] ^ DATA[7] ^ DATA[11] ^ DATA[19] ^ DATA[20] ^ DATA[21] ^ DATA[23] ^ DATA[24] ^ DATA[25] ^ DATA[26] ^ DATA[27] ^ DATA[29] ^ DATA[32] ^ DATA[39] ^ DATA[40] ^ DATA[42] ^ DATA[43] ^ DATA[45];
  assign CRC_OUT[28] = CRC_IN[4] ^ CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[14] ^ CRC_IN[17] ^ CRC_IN[24] ^ CRC_IN[25] ^ CRC_IN[27] ^ CRC_IN[28] ^ CRC_IN[30] ^ DATA[2] ^ DATA[5] ^ DATA[6] ^ DATA[8] ^ DATA[12] ^ DATA[20] ^ DATA[21] ^ DATA[22] ^ DATA[24] ^ DATA[25] ^ DATA[26] ^ DATA[27] ^ DATA[28] ^ DATA[30] ^ DATA[33] ^ DATA[40] ^ DATA[41] ^ DATA[43] ^ DATA[44] ^ DATA[46];
  assign CRC_OUT[29] = CRC_IN[5] ^ CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[9] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[15] ^ CRC_IN[18] ^ CRC_IN[25] ^ CRC_IN[26] ^ CRC_IN[28] ^ CRC_IN[29] ^ CRC_IN[31] ^ DATA[3] ^ DATA[6] ^ DATA[7] ^ DATA[9] ^ DATA[13] ^ DATA[21] ^ DATA[22] ^ DATA[23] ^ DATA[25] ^ DATA[26] ^ DATA[27] ^ DATA[28] ^ DATA[29] ^ DATA[31] ^ DATA[34] ^ DATA[41] ^ DATA[42] ^ DATA[44] ^ DATA[45] ^ DATA[47];
  assign CRC_OUT[30] = CRC_IN[6] ^ CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[10] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[16] ^ CRC_IN[19] ^ CRC_IN[26] ^ CRC_IN[27] ^ CRC_IN[29] ^ CRC_IN[30] ^ DATA[4] ^ DATA[7] ^ DATA[8] ^ DATA[10] ^ DATA[14] ^ DATA[22] ^ DATA[23] ^ DATA[24] ^ DATA[26] ^ DATA[27] ^ DATA[28] ^ DATA[29] ^ DATA[30] ^ DATA[32] ^ DATA[35] ^ DATA[42] ^ DATA[43] ^ DATA[45] ^ DATA[46];
  assign CRC_OUT[31] = CRC_IN[7] ^ CRC_IN[8] ^ CRC_IN[9] ^ CRC_IN[11] ^ CRC_IN[12] ^ CRC_IN[13] ^ CRC_IN[14] ^ CRC_IN[15] ^ CRC_IN[17] ^ CRC_IN[20] ^ CRC_IN[27] ^ CRC_IN[28] ^ CRC_IN[30] ^ CRC_IN[31] ^ DATA[5] ^ DATA[8] ^ DATA[9] ^ DATA[11] ^ DATA[15] ^ DATA[23] ^ DATA[24] ^ DATA[25] ^ DATA[27] ^ DATA[28] ^ DATA[29] ^ DATA[30] ^ DATA[31] ^ DATA[33] ^ DATA[36] ^ DATA[43] ^ DATA[44] ^ DATA[46] ^ DATA[47];
endmodule
